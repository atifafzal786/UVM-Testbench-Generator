// Minimal tb_pkg.sv (placeholder)
package tb_pkg;
  // typedefs and common definitions
endpackage
