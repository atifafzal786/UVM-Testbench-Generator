// Minimal interface.sv (placeholder)
interface dut_if();
  // signals
endinterface
